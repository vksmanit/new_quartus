-- megafunction wizard: %ALTFP_MULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_MULT 

-- ============================================================
-- File Name: fp_mult.vhd
-- Megafunction Name(s):
-- 			ALTFP_MULT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2017  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_mult CBX_AUTO_BLACKBOX="ALL" DEDICATED_MULTIPLIER_CIRCUITRY="YES" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone IV E" EXCEPTION_HANDLING="NO" PIPELINE=5 REDUCED_FUNCTIONALITY="NO" ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 aclr clock dataa datab result
--VERSION_BEGIN 17.1 cbx_alt_ded_mult_y 2017:10:19:05:46:40:SJ cbx_altbarrel_shift 2017:10:19:05:46:40:SJ cbx_altera_mult_add 2017:10:19:05:46:40:SJ cbx_altera_mult_add_rtl 2017:10:19:05:46:40:SJ cbx_altfp_mult 2017:10:19:05:46:40:SJ cbx_altmult_add 2017:10:19:05:46:40:SJ cbx_cycloneii 2017:10:19:05:46:40:SJ cbx_lpm_add_sub 2017:10:19:05:46:40:SJ cbx_lpm_compare 2017:10:19:05:46:40:SJ cbx_lpm_mult 2017:10:19:05:46:40:SJ cbx_mgl 2017:10:19:06:38:12:SJ cbx_nadder 2017:10:19:05:46:40:SJ cbx_padd 2017:10:19:05:46:40:SJ cbx_parallel_add 2017:10:19:05:46:40:SJ cbx_stratix 2017:10:19:05:46:40:SJ cbx_stratixii 2017:10:19:05:46:40:SJ cbx_util_mgl 2017:10:19:05:46:40:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 4 lpm_mult 1 reg 136 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fp_mult_altfp_mult_v9o IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END fp_mult_altfp_mult_v9o;

 ARCHITECTURE RTL OF fp_mult_altfp_mult_v9o IS

	 SIGNAL	 dataa_exp_all_one_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dataa_exp_all_one_ff_p1_w_lg_q296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dataa_exp_all_one_ff_p1_w_lg_q291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_exp_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dataa_man_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q290w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dataa_man_not_zero_ff_p1_w_lg_q290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 dataa_man_not_zero_ff_p2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_exp_all_one_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_datab_exp_all_one_ff_p1_w_lg_q294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_datab_exp_all_one_ff_p1_w_lg_q289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 datab_exp_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 datab_man_not_zero_ff_p1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q288w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_datab_man_not_zero_ff_p1_w_lg_q288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 datab_man_not_zero_ff_p2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_exp2_bias	:	STD_LOGIC_VECTOR(9 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_exp_bias	:	STD_LOGIC_VECTOR(9 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 delay_man_product_msb	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_delay_man_product_msb_w_lg_q392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_delay_man_product_msb_w_lg_q394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 delay_man_product_msb_p0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_add_p1	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_ff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_is_infinity_ff1_w_lg_q462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_input_is_infinity_ff1_w_lg_q464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 input_is_nan_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_is_nan_ff1_w_lg_q474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 input_not_zero_dffe_0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_not_zero_dffe_1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_not_zero_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_input_not_zero_ff1_w_lg_q461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 lsb_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_result_ff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_p	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_round_p2	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range399w400w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range396w397w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_lg_w_q_range391w398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range399w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range396w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_round_p2_w_q_range391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 round_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sticky_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_exp_add_adder_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_add_adder_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_add_adder_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_lg_w_result_range454w455w456w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_result_range454w455w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_lg_w_result_range429w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_result	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range454w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_adj_adder_w_result_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_dataa	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_exp_bias_subtr_result	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_dataa	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_datab	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_round_adder_result	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range302w303w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range299w300w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range298w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_lg_w_result_range298w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_dataa	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_datab	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_result	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range302w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range299w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_product2_mult_w_result_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w478w479w480w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w_lg_w478w479w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w_lg_w468w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w478w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_man_result_round_range475w476w477w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_man_result_round_range465w466w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_inf_num459w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range81w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range91w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range101w107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range111w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range121w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range131w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range141w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range84w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range94w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range104w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range114w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range124w129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range134w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range144w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_result_round_range475w476w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_result_round_range465w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range403w406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range407w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range410w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range413w415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range416w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range419w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_all_one_range422w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_inf463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_zero453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range450w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w468w469w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_inf_num459w460w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w468w469w470w471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_is_inf457w458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_is_inf457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range227w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range233w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range239w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range245w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range251w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range263w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range157w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range269w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range275w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range281w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range81w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range91w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range101w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range111w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range121w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range131w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range163w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range169w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range175w176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range181w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range199w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_dataa_range205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range214w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range224w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range230w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range236w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range242w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range248w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range254w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range260w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range266w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range272w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range278w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range284w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range84w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range94w95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range104w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range124w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range134w135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range166w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range172w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range178w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range184w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range190w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range196w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range202w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_datab_range208w209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range433w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range436w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range438w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range440w441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range442w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range444w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_result_exp_not_zero_range448w449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range306w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range337w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range340w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range343w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range346w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range349w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range352w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range355w357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range358w360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range361w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range364w366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range310w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range367w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range370w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range313w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range316w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range319w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range322w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range325w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range328w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range331w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_range334w336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bias :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  dataa_exp_all_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  dataa_exp_not_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  dataa_man_not_zero :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  datab_exp_all_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  datab_exp_not_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  datab_man_not_zero :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  exp_is_inf :	STD_LOGIC;
	 SIGNAL  exp_is_zero :	STD_LOGIC;
	 SIGNAL  expmod :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  inf_num :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  lsb_bit :	STD_LOGIC;
	 SIGNAL  man_result_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_shift_full :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  result_exp_all_one :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  result_exp_not_zero :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  round_bit :	STD_LOGIC;
	 SIGNAL  round_carry :	STD_LOGIC;
	 SIGNAL  sticky_bit :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_all_one_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_exp_not_zero_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dataa_man_not_zero_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_all_one_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_exp_not_zero_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_datab_man_not_zero_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_result_round_range475w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_w_man_result_round_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_shift_full_range379w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_all_one_range422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_result_exp_not_zero_range450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_range334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop0 : FOR i IN 0 TO 21 GENERATE 
		wire_w_lg_w_lg_w478w479w480w(i) <= wire_w_lg_w478w479w(i) AND wire_input_is_nan_ff1_w_lg_q474w(0);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 21 GENERATE 
		wire_w_lg_w478w479w(i) <= wire_w478w(i) AND wire_w_lg_exp_is_zero453w(0);
	END GENERATE loop1;
	wire_w_lg_w468w469w(0) <= wire_w468w(0) AND wire_w_lg_exp_is_zero453w(0);
	loop2 : FOR i IN 0 TO 21 GENERATE 
		wire_w478w(i) <= wire_w_lg_w_lg_w_man_result_round_range475w476w477w(i) AND wire_w_lg_exp_is_inf463w(0);
	END GENERATE loop2;
	wire_w468w(0) <= wire_w_lg_w_lg_w_man_result_round_range465w466w467w(0) AND wire_w_lg_exp_is_inf463w(0);
	loop3 : FOR i IN 0 TO 21 GENERATE 
		wire_w_lg_w_lg_w_man_result_round_range475w476w477w(i) <= wire_w_lg_w_man_result_round_range475w476w(i) AND wire_input_is_infinity_ff1_w_lg_q464w(0);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_man_result_round_range465w466w467w(0) <= wire_w_lg_w_man_result_round_range465w466w(0) AND wire_input_is_infinity_ff1_w_lg_q464w(0);
	loop4 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_inf_num459w(i) <= inf_num(i) AND wire_w_lg_w_lg_exp_is_inf457w458w(0);
	END GENERATE loop4;
	wire_w_lg_w_dataa_range81w87w(0) <= wire_w_dataa_range81w(0) AND wire_w_dataa_exp_all_one_range77w(0);
	wire_w_lg_w_dataa_range91w97w(0) <= wire_w_dataa_range91w(0) AND wire_w_dataa_exp_all_one_range88w(0);
	wire_w_lg_w_dataa_range101w107w(0) <= wire_w_dataa_range101w(0) AND wire_w_dataa_exp_all_one_range98w(0);
	wire_w_lg_w_dataa_range111w117w(0) <= wire_w_dataa_range111w(0) AND wire_w_dataa_exp_all_one_range108w(0);
	wire_w_lg_w_dataa_range121w127w(0) <= wire_w_dataa_range121w(0) AND wire_w_dataa_exp_all_one_range118w(0);
	wire_w_lg_w_dataa_range131w137w(0) <= wire_w_dataa_range131w(0) AND wire_w_dataa_exp_all_one_range128w(0);
	wire_w_lg_w_dataa_range141w147w(0) <= wire_w_dataa_range141w(0) AND wire_w_dataa_exp_all_one_range138w(0);
	wire_w_lg_w_datab_range84w89w(0) <= wire_w_datab_range84w(0) AND wire_w_datab_exp_all_one_range79w(0);
	wire_w_lg_w_datab_range94w99w(0) <= wire_w_datab_range94w(0) AND wire_w_datab_exp_all_one_range90w(0);
	wire_w_lg_w_datab_range104w109w(0) <= wire_w_datab_range104w(0) AND wire_w_datab_exp_all_one_range100w(0);
	wire_w_lg_w_datab_range114w119w(0) <= wire_w_datab_range114w(0) AND wire_w_datab_exp_all_one_range110w(0);
	wire_w_lg_w_datab_range124w129w(0) <= wire_w_datab_range124w(0) AND wire_w_datab_exp_all_one_range120w(0);
	wire_w_lg_w_datab_range134w139w(0) <= wire_w_datab_range134w(0) AND wire_w_datab_exp_all_one_range130w(0);
	wire_w_lg_w_datab_range144w149w(0) <= wire_w_datab_range144w(0) AND wire_w_datab_exp_all_one_range140w(0);
	loop5 : FOR i IN 0 TO 21 GENERATE 
		wire_w_lg_w_man_result_round_range475w476w(i) <= wire_w_man_result_round_range475w(i) AND input_not_zero_ff1;
	END GENERATE loop5;
	wire_w_lg_w_man_result_round_range465w466w(0) <= wire_w_man_result_round_range465w(0) AND input_not_zero_ff1;
	wire_w_lg_w_result_exp_all_one_range403w406w(0) <= wire_w_result_exp_all_one_range403w(0) AND wire_exp_adj_adder_w_result_range405w(0);
	wire_w_lg_w_result_exp_all_one_range407w409w(0) <= wire_w_result_exp_all_one_range407w(0) AND wire_exp_adj_adder_w_result_range408w(0);
	wire_w_lg_w_result_exp_all_one_range410w412w(0) <= wire_w_result_exp_all_one_range410w(0) AND wire_exp_adj_adder_w_result_range411w(0);
	wire_w_lg_w_result_exp_all_one_range413w415w(0) <= wire_w_result_exp_all_one_range413w(0) AND wire_exp_adj_adder_w_result_range414w(0);
	wire_w_lg_w_result_exp_all_one_range416w418w(0) <= wire_w_result_exp_all_one_range416w(0) AND wire_exp_adj_adder_w_result_range417w(0);
	wire_w_lg_w_result_exp_all_one_range419w421w(0) <= wire_w_result_exp_all_one_range419w(0) AND wire_exp_adj_adder_w_result_range420w(0);
	wire_w_lg_w_result_exp_all_one_range422w424w(0) <= wire_w_result_exp_all_one_range422w(0) AND wire_exp_adj_adder_w_result_range423w(0);
	wire_w_lg_exp_is_inf463w(0) <= NOT exp_is_inf;
	wire_w_lg_exp_is_zero453w(0) <= NOT exp_is_zero;
	wire_w_lg_w_result_exp_not_zero_range450w451w(0) <= NOT wire_w_result_exp_not_zero_range450w(0);
	wire_w_lg_w_lg_w468w469w470w(0) <= wire_w_lg_w468w469w(0) OR wire_input_is_infinity_ff1_w_lg_q462w(0);
	loop6 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_inf_num459w460w(i) <= wire_w_lg_inf_num459w(i) OR wire_exp_adj_adder_w_lg_w_lg_w_result_range454w455w456w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_w468w469w470w471w(0) <= wire_w_lg_w_lg_w468w469w470w(0) OR input_is_nan_ff1;
	wire_w_lg_w_lg_exp_is_inf457w458w(0) <= wire_w_lg_exp_is_inf457w(0) OR input_is_nan_ff1;
	wire_w_lg_exp_is_inf457w(0) <= exp_is_inf OR input_is_infinity_ff1;
	wire_w_lg_w_dataa_range211w212w(0) <= wire_w_dataa_range211w(0) OR wire_w_dataa_man_not_zero_range207w(0);
	wire_w_lg_w_dataa_range221w222w(0) <= wire_w_dataa_range221w(0) OR wire_w_dataa_man_not_zero_range218w(0);
	wire_w_lg_w_dataa_range227w228w(0) <= wire_w_dataa_range227w(0) OR wire_w_dataa_man_not_zero_range223w(0);
	wire_w_lg_w_dataa_range233w234w(0) <= wire_w_dataa_range233w(0) OR wire_w_dataa_man_not_zero_range229w(0);
	wire_w_lg_w_dataa_range239w240w(0) <= wire_w_dataa_range239w(0) OR wire_w_dataa_man_not_zero_range235w(0);
	wire_w_lg_w_dataa_range245w246w(0) <= wire_w_dataa_range245w(0) OR wire_w_dataa_man_not_zero_range241w(0);
	wire_w_lg_w_dataa_range251w252w(0) <= wire_w_dataa_range251w(0) OR wire_w_dataa_man_not_zero_range247w(0);
	wire_w_lg_w_dataa_range257w258w(0) <= wire_w_dataa_range257w(0) OR wire_w_dataa_man_not_zero_range253w(0);
	wire_w_lg_w_dataa_range263w264w(0) <= wire_w_dataa_range263w(0) OR wire_w_dataa_man_not_zero_range259w(0);
	wire_w_lg_w_dataa_range157w158w(0) <= wire_w_dataa_range157w(0) OR wire_w_dataa_man_not_zero_range152w(0);
	wire_w_lg_w_dataa_range269w270w(0) <= wire_w_dataa_range269w(0) OR wire_w_dataa_man_not_zero_range265w(0);
	wire_w_lg_w_dataa_range275w276w(0) <= wire_w_dataa_range275w(0) OR wire_w_dataa_man_not_zero_range271w(0);
	wire_w_lg_w_dataa_range281w282w(0) <= wire_w_dataa_range281w(0) OR wire_w_dataa_man_not_zero_range277w(0);
	wire_w_lg_w_dataa_range81w82w(0) <= wire_w_dataa_range81w(0) OR wire_w_dataa_exp_not_zero_range72w(0);
	wire_w_lg_w_dataa_range91w92w(0) <= wire_w_dataa_range91w(0) OR wire_w_dataa_exp_not_zero_range83w(0);
	wire_w_lg_w_dataa_range101w102w(0) <= wire_w_dataa_range101w(0) OR wire_w_dataa_exp_not_zero_range93w(0);
	wire_w_lg_w_dataa_range111w112w(0) <= wire_w_dataa_range111w(0) OR wire_w_dataa_exp_not_zero_range103w(0);
	wire_w_lg_w_dataa_range121w122w(0) <= wire_w_dataa_range121w(0) OR wire_w_dataa_exp_not_zero_range113w(0);
	wire_w_lg_w_dataa_range131w132w(0) <= wire_w_dataa_range131w(0) OR wire_w_dataa_exp_not_zero_range123w(0);
	wire_w_lg_w_dataa_range163w164w(0) <= wire_w_dataa_range163w(0) OR wire_w_dataa_man_not_zero_range159w(0);
	wire_w_lg_w_dataa_range141w142w(0) <= wire_w_dataa_range141w(0) OR wire_w_dataa_exp_not_zero_range133w(0);
	wire_w_lg_w_dataa_range169w170w(0) <= wire_w_dataa_range169w(0) OR wire_w_dataa_man_not_zero_range165w(0);
	wire_w_lg_w_dataa_range175w176w(0) <= wire_w_dataa_range175w(0) OR wire_w_dataa_man_not_zero_range171w(0);
	wire_w_lg_w_dataa_range181w182w(0) <= wire_w_dataa_range181w(0) OR wire_w_dataa_man_not_zero_range177w(0);
	wire_w_lg_w_dataa_range187w188w(0) <= wire_w_dataa_range187w(0) OR wire_w_dataa_man_not_zero_range183w(0);
	wire_w_lg_w_dataa_range193w194w(0) <= wire_w_dataa_range193w(0) OR wire_w_dataa_man_not_zero_range189w(0);
	wire_w_lg_w_dataa_range199w200w(0) <= wire_w_dataa_range199w(0) OR wire_w_dataa_man_not_zero_range195w(0);
	wire_w_lg_w_dataa_range205w206w(0) <= wire_w_dataa_range205w(0) OR wire_w_dataa_man_not_zero_range201w(0);
	wire_w_lg_w_datab_range214w215w(0) <= wire_w_datab_range214w(0) OR wire_w_datab_man_not_zero_range210w(0);
	wire_w_lg_w_datab_range224w225w(0) <= wire_w_datab_range224w(0) OR wire_w_datab_man_not_zero_range220w(0);
	wire_w_lg_w_datab_range230w231w(0) <= wire_w_datab_range230w(0) OR wire_w_datab_man_not_zero_range226w(0);
	wire_w_lg_w_datab_range236w237w(0) <= wire_w_datab_range236w(0) OR wire_w_datab_man_not_zero_range232w(0);
	wire_w_lg_w_datab_range242w243w(0) <= wire_w_datab_range242w(0) OR wire_w_datab_man_not_zero_range238w(0);
	wire_w_lg_w_datab_range248w249w(0) <= wire_w_datab_range248w(0) OR wire_w_datab_man_not_zero_range244w(0);
	wire_w_lg_w_datab_range254w255w(0) <= wire_w_datab_range254w(0) OR wire_w_datab_man_not_zero_range250w(0);
	wire_w_lg_w_datab_range260w261w(0) <= wire_w_datab_range260w(0) OR wire_w_datab_man_not_zero_range256w(0);
	wire_w_lg_w_datab_range266w267w(0) <= wire_w_datab_range266w(0) OR wire_w_datab_man_not_zero_range262w(0);
	wire_w_lg_w_datab_range160w161w(0) <= wire_w_datab_range160w(0) OR wire_w_datab_man_not_zero_range155w(0);
	wire_w_lg_w_datab_range272w273w(0) <= wire_w_datab_range272w(0) OR wire_w_datab_man_not_zero_range268w(0);
	wire_w_lg_w_datab_range278w279w(0) <= wire_w_datab_range278w(0) OR wire_w_datab_man_not_zero_range274w(0);
	wire_w_lg_w_datab_range284w285w(0) <= wire_w_datab_range284w(0) OR wire_w_datab_man_not_zero_range280w(0);
	wire_w_lg_w_datab_range84w85w(0) <= wire_w_datab_range84w(0) OR wire_w_datab_exp_not_zero_range75w(0);
	wire_w_lg_w_datab_range94w95w(0) <= wire_w_datab_range94w(0) OR wire_w_datab_exp_not_zero_range86w(0);
	wire_w_lg_w_datab_range104w105w(0) <= wire_w_datab_range104w(0) OR wire_w_datab_exp_not_zero_range96w(0);
	wire_w_lg_w_datab_range114w115w(0) <= wire_w_datab_range114w(0) OR wire_w_datab_exp_not_zero_range106w(0);
	wire_w_lg_w_datab_range124w125w(0) <= wire_w_datab_range124w(0) OR wire_w_datab_exp_not_zero_range116w(0);
	wire_w_lg_w_datab_range134w135w(0) <= wire_w_datab_range134w(0) OR wire_w_datab_exp_not_zero_range126w(0);
	wire_w_lg_w_datab_range166w167w(0) <= wire_w_datab_range166w(0) OR wire_w_datab_man_not_zero_range162w(0);
	wire_w_lg_w_datab_range144w145w(0) <= wire_w_datab_range144w(0) OR wire_w_datab_exp_not_zero_range136w(0);
	wire_w_lg_w_datab_range172w173w(0) <= wire_w_datab_range172w(0) OR wire_w_datab_man_not_zero_range168w(0);
	wire_w_lg_w_datab_range178w179w(0) <= wire_w_datab_range178w(0) OR wire_w_datab_man_not_zero_range174w(0);
	wire_w_lg_w_datab_range184w185w(0) <= wire_w_datab_range184w(0) OR wire_w_datab_man_not_zero_range180w(0);
	wire_w_lg_w_datab_range190w191w(0) <= wire_w_datab_range190w(0) OR wire_w_datab_man_not_zero_range186w(0);
	wire_w_lg_w_datab_range196w197w(0) <= wire_w_datab_range196w(0) OR wire_w_datab_man_not_zero_range192w(0);
	wire_w_lg_w_datab_range202w203w(0) <= wire_w_datab_range202w(0) OR wire_w_datab_man_not_zero_range198w(0);
	wire_w_lg_w_datab_range208w209w(0) <= wire_w_datab_range208w(0) OR wire_w_datab_man_not_zero_range204w(0);
	wire_w_lg_w_result_exp_not_zero_range433w435w(0) <= wire_w_result_exp_not_zero_range433w(0) OR wire_exp_adj_adder_w_result_range405w(0);
	wire_w_lg_w_result_exp_not_zero_range436w437w(0) <= wire_w_result_exp_not_zero_range436w(0) OR wire_exp_adj_adder_w_result_range408w(0);
	wire_w_lg_w_result_exp_not_zero_range438w439w(0) <= wire_w_result_exp_not_zero_range438w(0) OR wire_exp_adj_adder_w_result_range411w(0);
	wire_w_lg_w_result_exp_not_zero_range440w441w(0) <= wire_w_result_exp_not_zero_range440w(0) OR wire_exp_adj_adder_w_result_range414w(0);
	wire_w_lg_w_result_exp_not_zero_range442w443w(0) <= wire_w_result_exp_not_zero_range442w(0) OR wire_exp_adj_adder_w_result_range417w(0);
	wire_w_lg_w_result_exp_not_zero_range444w445w(0) <= wire_w_result_exp_not_zero_range444w(0) OR wire_exp_adj_adder_w_result_range420w(0);
	wire_w_lg_w_result_exp_not_zero_range446w447w(0) <= wire_w_result_exp_not_zero_range446w(0) OR wire_exp_adj_adder_w_result_range423w(0);
	wire_w_lg_w_result_exp_not_zero_range448w449w(0) <= wire_w_result_exp_not_zero_range448w(0) OR wire_exp_adj_adder_w_result_range426w(0);
	wire_w_lg_w_sticky_bit_range306w309w(0) <= wire_w_sticky_bit_range306w(0) OR wire_man_product2_mult_w_result_range308w(0);
	wire_w_lg_w_sticky_bit_range337w339w(0) <= wire_w_sticky_bit_range337w(0) OR wire_man_product2_mult_w_result_range338w(0);
	wire_w_lg_w_sticky_bit_range340w342w(0) <= wire_w_sticky_bit_range340w(0) OR wire_man_product2_mult_w_result_range341w(0);
	wire_w_lg_w_sticky_bit_range343w345w(0) <= wire_w_sticky_bit_range343w(0) OR wire_man_product2_mult_w_result_range344w(0);
	wire_w_lg_w_sticky_bit_range346w348w(0) <= wire_w_sticky_bit_range346w(0) OR wire_man_product2_mult_w_result_range347w(0);
	wire_w_lg_w_sticky_bit_range349w351w(0) <= wire_w_sticky_bit_range349w(0) OR wire_man_product2_mult_w_result_range350w(0);
	wire_w_lg_w_sticky_bit_range352w354w(0) <= wire_w_sticky_bit_range352w(0) OR wire_man_product2_mult_w_result_range353w(0);
	wire_w_lg_w_sticky_bit_range355w357w(0) <= wire_w_sticky_bit_range355w(0) OR wire_man_product2_mult_w_result_range356w(0);
	wire_w_lg_w_sticky_bit_range358w360w(0) <= wire_w_sticky_bit_range358w(0) OR wire_man_product2_mult_w_result_range359w(0);
	wire_w_lg_w_sticky_bit_range361w363w(0) <= wire_w_sticky_bit_range361w(0) OR wire_man_product2_mult_w_result_range362w(0);
	wire_w_lg_w_sticky_bit_range364w366w(0) <= wire_w_sticky_bit_range364w(0) OR wire_man_product2_mult_w_result_range365w(0);
	wire_w_lg_w_sticky_bit_range310w312w(0) <= wire_w_sticky_bit_range310w(0) OR wire_man_product2_mult_w_result_range311w(0);
	wire_w_lg_w_sticky_bit_range367w369w(0) <= wire_w_sticky_bit_range367w(0) OR wire_man_product2_mult_w_result_range368w(0);
	wire_w_lg_w_sticky_bit_range370w373w(0) <= wire_w_sticky_bit_range370w(0) OR wire_man_product2_mult_w_lg_w_result_range298w372w(0);
	wire_w_lg_w_sticky_bit_range313w315w(0) <= wire_w_sticky_bit_range313w(0) OR wire_man_product2_mult_w_result_range314w(0);
	wire_w_lg_w_sticky_bit_range316w318w(0) <= wire_w_sticky_bit_range316w(0) OR wire_man_product2_mult_w_result_range317w(0);
	wire_w_lg_w_sticky_bit_range319w321w(0) <= wire_w_sticky_bit_range319w(0) OR wire_man_product2_mult_w_result_range320w(0);
	wire_w_lg_w_sticky_bit_range322w324w(0) <= wire_w_sticky_bit_range322w(0) OR wire_man_product2_mult_w_result_range323w(0);
	wire_w_lg_w_sticky_bit_range325w327w(0) <= wire_w_sticky_bit_range325w(0) OR wire_man_product2_mult_w_result_range326w(0);
	wire_w_lg_w_sticky_bit_range328w330w(0) <= wire_w_sticky_bit_range328w(0) OR wire_man_product2_mult_w_result_range329w(0);
	wire_w_lg_w_sticky_bit_range331w333w(0) <= wire_w_sticky_bit_range331w(0) OR wire_man_product2_mult_w_result_range332w(0);
	wire_w_lg_w_sticky_bit_range334w336w(0) <= wire_w_sticky_bit_range334w(0) OR wire_man_product2_mult_w_result_range335w(0);
	bias <= ( "0" & "0" & "0" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	clk_en <= '1';
	dataa_exp_all_one <= ( wire_w_lg_w_dataa_range141w147w & wire_w_lg_w_dataa_range131w137w & wire_w_lg_w_dataa_range121w127w & wire_w_lg_w_dataa_range111w117w & wire_w_lg_w_dataa_range101w107w & wire_w_lg_w_dataa_range91w97w & wire_w_lg_w_dataa_range81w87w & dataa(23));
	dataa_exp_not_zero <= ( wire_w_lg_w_dataa_range141w142w & wire_w_lg_w_dataa_range131w132w & wire_w_lg_w_dataa_range121w122w & wire_w_lg_w_dataa_range111w112w & wire_w_lg_w_dataa_range101w102w & wire_w_lg_w_dataa_range91w92w & wire_w_lg_w_dataa_range81w82w & dataa(23));
	dataa_man_not_zero <= ( wire_w_lg_w_dataa_range281w282w & wire_w_lg_w_dataa_range275w276w & wire_w_lg_w_dataa_range269w270w & wire_w_lg_w_dataa_range263w264w & wire_w_lg_w_dataa_range257w258w & wire_w_lg_w_dataa_range251w252w & wire_w_lg_w_dataa_range245w246w & wire_w_lg_w_dataa_range239w240w & wire_w_lg_w_dataa_range233w234w & wire_w_lg_w_dataa_range227w228w & wire_w_lg_w_dataa_range221w222w & dataa(11) & wire_w_lg_w_dataa_range211w212w & wire_w_lg_w_dataa_range205w206w & wire_w_lg_w_dataa_range199w200w & wire_w_lg_w_dataa_range193w194w & wire_w_lg_w_dataa_range187w188w & wire_w_lg_w_dataa_range181w182w & wire_w_lg_w_dataa_range175w176w & wire_w_lg_w_dataa_range169w170w & wire_w_lg_w_dataa_range163w164w & wire_w_lg_w_dataa_range157w158w & dataa(0));
	datab_exp_all_one <= ( wire_w_lg_w_datab_range144w149w & wire_w_lg_w_datab_range134w139w & wire_w_lg_w_datab_range124w129w & wire_w_lg_w_datab_range114w119w & wire_w_lg_w_datab_range104w109w & wire_w_lg_w_datab_range94w99w & wire_w_lg_w_datab_range84w89w & datab(23));
	datab_exp_not_zero <= ( wire_w_lg_w_datab_range144w145w & wire_w_lg_w_datab_range134w135w & wire_w_lg_w_datab_range124w125w & wire_w_lg_w_datab_range114w115w & wire_w_lg_w_datab_range104w105w & wire_w_lg_w_datab_range94w95w & wire_w_lg_w_datab_range84w85w & datab(23));
	datab_man_not_zero <= ( wire_w_lg_w_datab_range284w285w & wire_w_lg_w_datab_range278w279w & wire_w_lg_w_datab_range272w273w & wire_w_lg_w_datab_range266w267w & wire_w_lg_w_datab_range260w261w & wire_w_lg_w_datab_range254w255w & wire_w_lg_w_datab_range248w249w & wire_w_lg_w_datab_range242w243w & wire_w_lg_w_datab_range236w237w & wire_w_lg_w_datab_range230w231w & wire_w_lg_w_datab_range224w225w & datab(11) & wire_w_lg_w_datab_range214w215w & wire_w_lg_w_datab_range208w209w & wire_w_lg_w_datab_range202w203w & wire_w_lg_w_datab_range196w197w & wire_w_lg_w_datab_range190w191w & wire_w_lg_w_datab_range184w185w & wire_w_lg_w_datab_range178w179w & wire_w_lg_w_datab_range172w173w & wire_w_lg_w_datab_range166w167w & wire_w_lg_w_datab_range160w161w & datab(0));
	exp_is_inf <= (((NOT wire_exp_adj_adder_result(9)) AND wire_exp_adj_adder_result(8)) OR ((NOT wire_exp_adj_adder_result(8)) AND result_exp_all_one(7)));
	exp_is_zero <= wire_exp_adj_adder_w_lg_w_result_range429w452w(0);
	expmod <= ( "00000000" & wire_delay_man_product_msb_w_lg_q392w & wire_delay_man_product_msb_w_lg_q394w);
	inf_num <= ( "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	lsb_bit <= man_shift_full(1);
	man_result_round <= (wire_man_round_p2_w_lg_w_q_range399w400w OR wire_man_round_p2_w_lg_w_q_range396w397w);
	man_shift_full <= (wire_man_product2_mult_w_lg_w_result_range302w303w OR wire_man_product2_mult_w_lg_w_result_range299w300w);
	result <= ( sign_node_ff4 & exp_result_ff(7 DOWNTO 0) & man_result_ff(22 DOWNTO 0));
	result_exp_all_one <= ( wire_w_lg_w_result_exp_all_one_range422w424w & wire_w_lg_w_result_exp_all_one_range419w421w & wire_w_lg_w_result_exp_all_one_range416w418w & wire_w_lg_w_result_exp_all_one_range413w415w & wire_w_lg_w_result_exp_all_one_range410w412w & wire_w_lg_w_result_exp_all_one_range407w409w & wire_w_lg_w_result_exp_all_one_range403w406w & wire_exp_adj_adder_result(0));
	result_exp_not_zero <= ( wire_w_lg_w_result_exp_not_zero_range448w449w & wire_w_lg_w_result_exp_not_zero_range446w447w & wire_w_lg_w_result_exp_not_zero_range444w445w & wire_w_lg_w_result_exp_not_zero_range442w443w & wire_w_lg_w_result_exp_not_zero_range440w441w & wire_w_lg_w_result_exp_not_zero_range438w439w & wire_w_lg_w_result_exp_not_zero_range436w437w & wire_w_lg_w_result_exp_not_zero_range433w435w & wire_exp_adj_adder_result(0));
	round_bit <= man_shift_full(0);
	round_carry <= (round_dffe AND (lsb_dffe OR sticky_dffe));
	sticky_bit <= ( wire_w_lg_w_sticky_bit_range370w373w & wire_w_lg_w_sticky_bit_range367w369w & wire_w_lg_w_sticky_bit_range364w366w & wire_w_lg_w_sticky_bit_range361w363w & wire_w_lg_w_sticky_bit_range358w360w & wire_w_lg_w_sticky_bit_range355w357w & wire_w_lg_w_sticky_bit_range352w354w & wire_w_lg_w_sticky_bit_range349w351w & wire_w_lg_w_sticky_bit_range346w348w & wire_w_lg_w_sticky_bit_range343w345w & wire_w_lg_w_sticky_bit_range340w342w & wire_w_lg_w_sticky_bit_range337w339w & wire_w_lg_w_sticky_bit_range334w336w & wire_w_lg_w_sticky_bit_range331w333w & wire_w_lg_w_sticky_bit_range328w330w & wire_w_lg_w_sticky_bit_range325w327w & wire_w_lg_w_sticky_bit_range322w324w & wire_w_lg_w_sticky_bit_range319w321w & wire_w_lg_w_sticky_bit_range316w318w & wire_w_lg_w_sticky_bit_range313w315w & wire_w_lg_w_sticky_bit_range310w312w & wire_w_lg_w_sticky_bit_range306w309w & wire_man_product2_mult_result(0));
	wire_w_dataa_range211w(0) <= dataa(10);
	wire_w_dataa_range221w(0) <= dataa(12);
	wire_w_dataa_range227w(0) <= dataa(13);
	wire_w_dataa_range233w(0) <= dataa(14);
	wire_w_dataa_range239w(0) <= dataa(15);
	wire_w_dataa_range245w(0) <= dataa(16);
	wire_w_dataa_range251w(0) <= dataa(17);
	wire_w_dataa_range257w(0) <= dataa(18);
	wire_w_dataa_range263w(0) <= dataa(19);
	wire_w_dataa_range157w(0) <= dataa(1);
	wire_w_dataa_range269w(0) <= dataa(20);
	wire_w_dataa_range275w(0) <= dataa(21);
	wire_w_dataa_range281w(0) <= dataa(22);
	wire_w_dataa_range81w(0) <= dataa(24);
	wire_w_dataa_range91w(0) <= dataa(25);
	wire_w_dataa_range101w(0) <= dataa(26);
	wire_w_dataa_range111w(0) <= dataa(27);
	wire_w_dataa_range121w(0) <= dataa(28);
	wire_w_dataa_range131w(0) <= dataa(29);
	wire_w_dataa_range163w(0) <= dataa(2);
	wire_w_dataa_range141w(0) <= dataa(30);
	wire_w_dataa_range169w(0) <= dataa(3);
	wire_w_dataa_range175w(0) <= dataa(4);
	wire_w_dataa_range181w(0) <= dataa(5);
	wire_w_dataa_range187w(0) <= dataa(6);
	wire_w_dataa_range193w(0) <= dataa(7);
	wire_w_dataa_range199w(0) <= dataa(8);
	wire_w_dataa_range205w(0) <= dataa(9);
	wire_w_dataa_exp_all_one_range77w(0) <= dataa_exp_all_one(0);
	wire_w_dataa_exp_all_one_range88w(0) <= dataa_exp_all_one(1);
	wire_w_dataa_exp_all_one_range98w(0) <= dataa_exp_all_one(2);
	wire_w_dataa_exp_all_one_range108w(0) <= dataa_exp_all_one(3);
	wire_w_dataa_exp_all_one_range118w(0) <= dataa_exp_all_one(4);
	wire_w_dataa_exp_all_one_range128w(0) <= dataa_exp_all_one(5);
	wire_w_dataa_exp_all_one_range138w(0) <= dataa_exp_all_one(6);
	wire_w_dataa_exp_not_zero_range72w(0) <= dataa_exp_not_zero(0);
	wire_w_dataa_exp_not_zero_range83w(0) <= dataa_exp_not_zero(1);
	wire_w_dataa_exp_not_zero_range93w(0) <= dataa_exp_not_zero(2);
	wire_w_dataa_exp_not_zero_range103w(0) <= dataa_exp_not_zero(3);
	wire_w_dataa_exp_not_zero_range113w(0) <= dataa_exp_not_zero(4);
	wire_w_dataa_exp_not_zero_range123w(0) <= dataa_exp_not_zero(5);
	wire_w_dataa_exp_not_zero_range133w(0) <= dataa_exp_not_zero(6);
	wire_w_dataa_man_not_zero_range152w(0) <= dataa_man_not_zero(0);
	wire_w_dataa_man_not_zero_range218w(0) <= dataa_man_not_zero(11);
	wire_w_dataa_man_not_zero_range223w(0) <= dataa_man_not_zero(12);
	wire_w_dataa_man_not_zero_range229w(0) <= dataa_man_not_zero(13);
	wire_w_dataa_man_not_zero_range235w(0) <= dataa_man_not_zero(14);
	wire_w_dataa_man_not_zero_range241w(0) <= dataa_man_not_zero(15);
	wire_w_dataa_man_not_zero_range247w(0) <= dataa_man_not_zero(16);
	wire_w_dataa_man_not_zero_range253w(0) <= dataa_man_not_zero(17);
	wire_w_dataa_man_not_zero_range259w(0) <= dataa_man_not_zero(18);
	wire_w_dataa_man_not_zero_range265w(0) <= dataa_man_not_zero(19);
	wire_w_dataa_man_not_zero_range159w(0) <= dataa_man_not_zero(1);
	wire_w_dataa_man_not_zero_range271w(0) <= dataa_man_not_zero(20);
	wire_w_dataa_man_not_zero_range277w(0) <= dataa_man_not_zero(21);
	wire_w_dataa_man_not_zero_range165w(0) <= dataa_man_not_zero(2);
	wire_w_dataa_man_not_zero_range171w(0) <= dataa_man_not_zero(3);
	wire_w_dataa_man_not_zero_range177w(0) <= dataa_man_not_zero(4);
	wire_w_dataa_man_not_zero_range183w(0) <= dataa_man_not_zero(5);
	wire_w_dataa_man_not_zero_range189w(0) <= dataa_man_not_zero(6);
	wire_w_dataa_man_not_zero_range195w(0) <= dataa_man_not_zero(7);
	wire_w_dataa_man_not_zero_range201w(0) <= dataa_man_not_zero(8);
	wire_w_dataa_man_not_zero_range207w(0) <= dataa_man_not_zero(9);
	wire_w_datab_range214w(0) <= datab(10);
	wire_w_datab_range224w(0) <= datab(12);
	wire_w_datab_range230w(0) <= datab(13);
	wire_w_datab_range236w(0) <= datab(14);
	wire_w_datab_range242w(0) <= datab(15);
	wire_w_datab_range248w(0) <= datab(16);
	wire_w_datab_range254w(0) <= datab(17);
	wire_w_datab_range260w(0) <= datab(18);
	wire_w_datab_range266w(0) <= datab(19);
	wire_w_datab_range160w(0) <= datab(1);
	wire_w_datab_range272w(0) <= datab(20);
	wire_w_datab_range278w(0) <= datab(21);
	wire_w_datab_range284w(0) <= datab(22);
	wire_w_datab_range84w(0) <= datab(24);
	wire_w_datab_range94w(0) <= datab(25);
	wire_w_datab_range104w(0) <= datab(26);
	wire_w_datab_range114w(0) <= datab(27);
	wire_w_datab_range124w(0) <= datab(28);
	wire_w_datab_range134w(0) <= datab(29);
	wire_w_datab_range166w(0) <= datab(2);
	wire_w_datab_range144w(0) <= datab(30);
	wire_w_datab_range172w(0) <= datab(3);
	wire_w_datab_range178w(0) <= datab(4);
	wire_w_datab_range184w(0) <= datab(5);
	wire_w_datab_range190w(0) <= datab(6);
	wire_w_datab_range196w(0) <= datab(7);
	wire_w_datab_range202w(0) <= datab(8);
	wire_w_datab_range208w(0) <= datab(9);
	wire_w_datab_exp_all_one_range79w(0) <= datab_exp_all_one(0);
	wire_w_datab_exp_all_one_range90w(0) <= datab_exp_all_one(1);
	wire_w_datab_exp_all_one_range100w(0) <= datab_exp_all_one(2);
	wire_w_datab_exp_all_one_range110w(0) <= datab_exp_all_one(3);
	wire_w_datab_exp_all_one_range120w(0) <= datab_exp_all_one(4);
	wire_w_datab_exp_all_one_range130w(0) <= datab_exp_all_one(5);
	wire_w_datab_exp_all_one_range140w(0) <= datab_exp_all_one(6);
	wire_w_datab_exp_not_zero_range75w(0) <= datab_exp_not_zero(0);
	wire_w_datab_exp_not_zero_range86w(0) <= datab_exp_not_zero(1);
	wire_w_datab_exp_not_zero_range96w(0) <= datab_exp_not_zero(2);
	wire_w_datab_exp_not_zero_range106w(0) <= datab_exp_not_zero(3);
	wire_w_datab_exp_not_zero_range116w(0) <= datab_exp_not_zero(4);
	wire_w_datab_exp_not_zero_range126w(0) <= datab_exp_not_zero(5);
	wire_w_datab_exp_not_zero_range136w(0) <= datab_exp_not_zero(6);
	wire_w_datab_man_not_zero_range155w(0) <= datab_man_not_zero(0);
	wire_w_datab_man_not_zero_range220w(0) <= datab_man_not_zero(11);
	wire_w_datab_man_not_zero_range226w(0) <= datab_man_not_zero(12);
	wire_w_datab_man_not_zero_range232w(0) <= datab_man_not_zero(13);
	wire_w_datab_man_not_zero_range238w(0) <= datab_man_not_zero(14);
	wire_w_datab_man_not_zero_range244w(0) <= datab_man_not_zero(15);
	wire_w_datab_man_not_zero_range250w(0) <= datab_man_not_zero(16);
	wire_w_datab_man_not_zero_range256w(0) <= datab_man_not_zero(17);
	wire_w_datab_man_not_zero_range262w(0) <= datab_man_not_zero(18);
	wire_w_datab_man_not_zero_range268w(0) <= datab_man_not_zero(19);
	wire_w_datab_man_not_zero_range162w(0) <= datab_man_not_zero(1);
	wire_w_datab_man_not_zero_range274w(0) <= datab_man_not_zero(20);
	wire_w_datab_man_not_zero_range280w(0) <= datab_man_not_zero(21);
	wire_w_datab_man_not_zero_range168w(0) <= datab_man_not_zero(2);
	wire_w_datab_man_not_zero_range174w(0) <= datab_man_not_zero(3);
	wire_w_datab_man_not_zero_range180w(0) <= datab_man_not_zero(4);
	wire_w_datab_man_not_zero_range186w(0) <= datab_man_not_zero(5);
	wire_w_datab_man_not_zero_range192w(0) <= datab_man_not_zero(6);
	wire_w_datab_man_not_zero_range198w(0) <= datab_man_not_zero(7);
	wire_w_datab_man_not_zero_range204w(0) <= datab_man_not_zero(8);
	wire_w_datab_man_not_zero_range210w(0) <= datab_man_not_zero(9);
	wire_w_man_result_round_range475w <= man_result_round(21 DOWNTO 0);
	wire_w_man_result_round_range465w(0) <= man_result_round(22);
	wire_w_man_shift_full_range379w <= man_shift_full(24 DOWNTO 1);
	wire_w_result_exp_all_one_range403w(0) <= result_exp_all_one(0);
	wire_w_result_exp_all_one_range407w(0) <= result_exp_all_one(1);
	wire_w_result_exp_all_one_range410w(0) <= result_exp_all_one(2);
	wire_w_result_exp_all_one_range413w(0) <= result_exp_all_one(3);
	wire_w_result_exp_all_one_range416w(0) <= result_exp_all_one(4);
	wire_w_result_exp_all_one_range419w(0) <= result_exp_all_one(5);
	wire_w_result_exp_all_one_range422w(0) <= result_exp_all_one(6);
	wire_w_result_exp_not_zero_range433w(0) <= result_exp_not_zero(0);
	wire_w_result_exp_not_zero_range436w(0) <= result_exp_not_zero(1);
	wire_w_result_exp_not_zero_range438w(0) <= result_exp_not_zero(2);
	wire_w_result_exp_not_zero_range440w(0) <= result_exp_not_zero(3);
	wire_w_result_exp_not_zero_range442w(0) <= result_exp_not_zero(4);
	wire_w_result_exp_not_zero_range444w(0) <= result_exp_not_zero(5);
	wire_w_result_exp_not_zero_range446w(0) <= result_exp_not_zero(6);
	wire_w_result_exp_not_zero_range448w(0) <= result_exp_not_zero(7);
	wire_w_result_exp_not_zero_range450w(0) <= result_exp_not_zero(8);
	wire_w_sticky_bit_range306w(0) <= sticky_bit(0);
	wire_w_sticky_bit_range337w(0) <= sticky_bit(10);
	wire_w_sticky_bit_range340w(0) <= sticky_bit(11);
	wire_w_sticky_bit_range343w(0) <= sticky_bit(12);
	wire_w_sticky_bit_range346w(0) <= sticky_bit(13);
	wire_w_sticky_bit_range349w(0) <= sticky_bit(14);
	wire_w_sticky_bit_range352w(0) <= sticky_bit(15);
	wire_w_sticky_bit_range355w(0) <= sticky_bit(16);
	wire_w_sticky_bit_range358w(0) <= sticky_bit(17);
	wire_w_sticky_bit_range361w(0) <= sticky_bit(18);
	wire_w_sticky_bit_range364w(0) <= sticky_bit(19);
	wire_w_sticky_bit_range310w(0) <= sticky_bit(1);
	wire_w_sticky_bit_range367w(0) <= sticky_bit(20);
	wire_w_sticky_bit_range370w(0) <= sticky_bit(21);
	wire_w_sticky_bit_range313w(0) <= sticky_bit(2);
	wire_w_sticky_bit_range316w(0) <= sticky_bit(3);
	wire_w_sticky_bit_range319w(0) <= sticky_bit(4);
	wire_w_sticky_bit_range322w(0) <= sticky_bit(5);
	wire_w_sticky_bit_range325w(0) <= sticky_bit(6);
	wire_w_sticky_bit_range328w(0) <= sticky_bit(7);
	wire_w_sticky_bit_range331w(0) <= sticky_bit(8);
	wire_w_sticky_bit_range334w(0) <= sticky_bit(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_exp_all_one_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_exp_all_one_ff_p1 <= dataa_exp_all_one(7);
			END IF;
		END IF;
	END PROCESS;
	wire_dataa_exp_all_one_ff_p1_w_lg_q296w(0) <= dataa_exp_all_one_ff_p1 AND wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q290w295w(0);
	wire_dataa_exp_all_one_ff_p1_w_lg_q291w(0) <= dataa_exp_all_one_ff_p1 AND wire_dataa_man_not_zero_ff_p1_w_lg_q290w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_exp_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_exp_not_zero_ff_p1 <= dataa_exp_not_zero(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_man_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_man_not_zero_ff_p1 <= dataa_man_not_zero(10);
			END IF;
		END IF;
	END PROCESS;
	wire_dataa_man_not_zero_ff_p1_w_lg_w_lg_q290w295w(0) <= NOT wire_dataa_man_not_zero_ff_p1_w_lg_q290w(0);
	wire_dataa_man_not_zero_ff_p1_w_lg_q290w(0) <= dataa_man_not_zero_ff_p1 OR dataa_man_not_zero_ff_p2;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dataa_man_not_zero_ff_p2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dataa_man_not_zero_ff_p2 <= dataa_man_not_zero(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_exp_all_one_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_exp_all_one_ff_p1 <= datab_exp_all_one(7);
			END IF;
		END IF;
	END PROCESS;
	wire_datab_exp_all_one_ff_p1_w_lg_q294w(0) <= datab_exp_all_one_ff_p1 AND wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q288w293w(0);
	wire_datab_exp_all_one_ff_p1_w_lg_q289w(0) <= datab_exp_all_one_ff_p1 AND wire_datab_man_not_zero_ff_p1_w_lg_q288w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_exp_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_exp_not_zero_ff_p1 <= datab_exp_not_zero(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_man_not_zero_ff_p1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_man_not_zero_ff_p1 <= datab_man_not_zero(10);
			END IF;
		END IF;
	END PROCESS;
	wire_datab_man_not_zero_ff_p1_w_lg_w_lg_q288w293w(0) <= NOT wire_datab_man_not_zero_ff_p1_w_lg_q288w(0);
	wire_datab_man_not_zero_ff_p1_w_lg_q288w(0) <= datab_man_not_zero_ff_p1 OR datab_man_not_zero_ff_p2;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN datab_man_not_zero_ff_p2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN datab_man_not_zero_ff_p2 <= datab_man_not_zero(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_exp2_bias <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_exp2_bias <= delay_exp_bias;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_exp_bias <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_exp_bias <= wire_exp_bias_subtr_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_man_product_msb <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_man_product_msb <= delay_man_product_msb_p0;
			END IF;
		END IF;
	END PROCESS;
	wire_delay_man_product_msb_w_lg_q392w(0) <= delay_man_product_msb AND wire_man_round_p2_w_q_range391w(0);
	wire_delay_man_product_msb_w_lg_q394w(0) <= delay_man_product_msb XOR wire_man_round_p2_w_q_range391w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN delay_man_product_msb_p0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN delay_man_product_msb_p0 <= wire_man_product2_mult_w_result_range298w(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_add_p1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_add_p1 <= wire_exp_add_adder_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_ff <= wire_w_lg_w_lg_inf_num459w460w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_dffe_0 <= (wire_dataa_exp_all_one_ff_p1_w_lg_q296w(0) OR wire_datab_exp_all_one_ff_p1_w_lg_q294w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_dffe_1 <= input_is_infinity_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_ff1 <= input_is_infinity_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_is_infinity_ff1_w_lg_q462w(0) <= input_is_infinity_ff1 AND wire_input_not_zero_ff1_w_lg_q461w(0);
	wire_input_is_infinity_ff1_w_lg_q464w(0) <= NOT input_is_infinity_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe_0 <= (wire_dataa_exp_all_one_ff_p1_w_lg_q291w(0) OR wire_datab_exp_all_one_ff_p1_w_lg_q289w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_dffe_1 <= input_is_nan_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_ff1 <= input_is_nan_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_is_nan_ff1_w_lg_q474w(0) <= NOT input_is_nan_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_dffe_0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_dffe_0 <= (dataa_exp_not_zero_ff_p1 AND datab_exp_not_zero_ff_p1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_dffe_1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_dffe_1 <= input_not_zero_dffe_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_not_zero_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_not_zero_ff1 <= input_not_zero_dffe_1;
			END IF;
		END IF;
	END PROCESS;
	wire_input_not_zero_ff1_w_lg_q461w(0) <= NOT input_not_zero_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lsb_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lsb_dffe <= lsb_bit;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_ff <= ( wire_w_lg_w_lg_w_lg_w468w469w470w471w & wire_w_lg_w_lg_w478w479w480w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_p <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_p <= wire_w_man_shift_full_range379w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_round_p2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_round_p2 <= wire_man_round_adder_result;
			END IF;
		END IF;
	END PROCESS;
	loop7 : FOR i IN 0 TO 23 GENERATE 
		wire_man_round_p2_w_lg_w_q_range399w400w(i) <= wire_man_round_p2_w_q_range399w(i) AND wire_man_round_p2_w_lg_w_q_range391w398w(0);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 23 GENERATE 
		wire_man_round_p2_w_lg_w_q_range396w397w(i) <= wire_man_round_p2_w_q_range396w(i) AND wire_man_round_p2_w_q_range391w(0);
	END GENERATE loop8;
	wire_man_round_p2_w_lg_w_q_range391w398w(0) <= NOT wire_man_round_p2_w_q_range391w(0);
	wire_man_round_p2_w_q_range399w <= man_round_p2(23 DOWNTO 0);
	wire_man_round_p2_w_q_range396w <= man_round_p2(24 DOWNTO 1);
	wire_man_round_p2_w_q_range391w(0) <= man_round_p2(24);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN round_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN round_dffe <= round_bit;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff0 <= (dataa(31) XOR datab(31));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff1 <= sign_node_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff2 <= sign_node_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff3 <= sign_node_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff4 <= sign_node_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sticky_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sticky_dffe <= sticky_bit(22);
			END IF;
		END IF;
	END PROCESS;
	wire_exp_add_adder_dataa <= ( "0" & dataa(30 DOWNTO 23));
	wire_exp_add_adder_datab <= ( "0" & datab(30 DOWNTO 23));
	exp_add_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clk_en,
		clock => clock,
		dataa => wire_exp_add_adder_dataa,
		datab => wire_exp_add_adder_datab,
		result => wire_exp_add_adder_result
	  );
	loop9 : FOR i IN 0 TO 7 GENERATE 
		wire_exp_adj_adder_w_lg_w_lg_w_result_range454w455w456w(i) <= wire_exp_adj_adder_w_lg_w_result_range454w455w(i) AND input_not_zero_ff1;
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 7 GENERATE 
		wire_exp_adj_adder_w_lg_w_result_range454w455w(i) <= wire_exp_adj_adder_w_result_range454w(i) AND wire_w_lg_exp_is_zero453w(0);
	END GENERATE loop10;
	wire_exp_adj_adder_w_lg_w_result_range429w452w(0) <= wire_exp_adj_adder_w_result_range429w(0) OR wire_w_lg_w_result_exp_not_zero_range450w451w(0);
	wire_exp_adj_adder_w_result_range405w(0) <= wire_exp_adj_adder_result(1);
	wire_exp_adj_adder_w_result_range408w(0) <= wire_exp_adj_adder_result(2);
	wire_exp_adj_adder_w_result_range411w(0) <= wire_exp_adj_adder_result(3);
	wire_exp_adj_adder_w_result_range414w(0) <= wire_exp_adj_adder_result(4);
	wire_exp_adj_adder_w_result_range417w(0) <= wire_exp_adj_adder_result(5);
	wire_exp_adj_adder_w_result_range420w(0) <= wire_exp_adj_adder_result(6);
	wire_exp_adj_adder_w_result_range454w <= wire_exp_adj_adder_result(7 DOWNTO 0);
	wire_exp_adj_adder_w_result_range423w(0) <= wire_exp_adj_adder_result(7);
	wire_exp_adj_adder_w_result_range426w(0) <= wire_exp_adj_adder_result(8);
	wire_exp_adj_adder_w_result_range429w(0) <= wire_exp_adj_adder_result(9);
	exp_adj_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 10
	  )
	  PORT MAP ( 
		cin => wire_gnd,
		dataa => delay_exp2_bias,
		datab => expmod,
		result => wire_exp_adj_adder_result
	  );
	wire_exp_bias_subtr_dataa <= ( "0" & exp_add_p1(8 DOWNTO 0));
	wire_exp_bias_subtr_datab <= ( bias(9 DOWNTO 0));
	exp_bias_subtr :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 0,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 10
	  )
	  PORT MAP ( 
		dataa => wire_exp_bias_subtr_dataa,
		datab => wire_exp_bias_subtr_datab,
		result => wire_exp_bias_subtr_result
	  );
	wire_man_round_adder_dataa <= ( "0" & man_round_p);
	wire_man_round_adder_datab <= ( "000000000000000000000000" & round_carry);
	man_round_adder :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 0,
		LPM_WIDTH => 25
	  )
	  PORT MAP ( 
		dataa => wire_man_round_adder_dataa,
		datab => wire_man_round_adder_datab,
		result => wire_man_round_adder_result
	  );
	loop11 : FOR i IN 0 TO 24 GENERATE 
		wire_man_product2_mult_w_lg_w_result_range302w303w(i) <= wire_man_product2_mult_w_result_range302w(i) AND wire_man_product2_mult_w_lg_w_result_range298w301w(0);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 24 GENERATE 
		wire_man_product2_mult_w_lg_w_result_range299w300w(i) <= wire_man_product2_mult_w_result_range299w(i) AND wire_man_product2_mult_w_result_range298w(0);
	END GENERATE loop12;
	wire_man_product2_mult_w_lg_w_result_range298w372w(0) <= wire_man_product2_mult_w_result_range298w(0) AND wire_man_product2_mult_w_result_range371w(0);
	wire_man_product2_mult_w_lg_w_result_range298w301w(0) <= NOT wire_man_product2_mult_w_result_range298w(0);
	wire_man_product2_mult_dataa <= ( "1" & dataa(22 DOWNTO 0));
	wire_man_product2_mult_datab <= ( "1" & datab(22 DOWNTO 0));
	wire_man_product2_mult_w_result_range335w(0) <= wire_man_product2_mult_result(10);
	wire_man_product2_mult_w_result_range338w(0) <= wire_man_product2_mult_result(11);
	wire_man_product2_mult_w_result_range341w(0) <= wire_man_product2_mult_result(12);
	wire_man_product2_mult_w_result_range344w(0) <= wire_man_product2_mult_result(13);
	wire_man_product2_mult_w_result_range347w(0) <= wire_man_product2_mult_result(14);
	wire_man_product2_mult_w_result_range350w(0) <= wire_man_product2_mult_result(15);
	wire_man_product2_mult_w_result_range353w(0) <= wire_man_product2_mult_result(16);
	wire_man_product2_mult_w_result_range356w(0) <= wire_man_product2_mult_result(17);
	wire_man_product2_mult_w_result_range359w(0) <= wire_man_product2_mult_result(18);
	wire_man_product2_mult_w_result_range362w(0) <= wire_man_product2_mult_result(19);
	wire_man_product2_mult_w_result_range308w(0) <= wire_man_product2_mult_result(1);
	wire_man_product2_mult_w_result_range365w(0) <= wire_man_product2_mult_result(20);
	wire_man_product2_mult_w_result_range368w(0) <= wire_man_product2_mult_result(21);
	wire_man_product2_mult_w_result_range371w(0) <= wire_man_product2_mult_result(22);
	wire_man_product2_mult_w_result_range311w(0) <= wire_man_product2_mult_result(2);
	wire_man_product2_mult_w_result_range314w(0) <= wire_man_product2_mult_result(3);
	wire_man_product2_mult_w_result_range302w <= wire_man_product2_mult_result(46 DOWNTO 22);
	wire_man_product2_mult_w_result_range299w <= wire_man_product2_mult_result(47 DOWNTO 23);
	wire_man_product2_mult_w_result_range298w(0) <= wire_man_product2_mult_result(47);
	wire_man_product2_mult_w_result_range317w(0) <= wire_man_product2_mult_result(4);
	wire_man_product2_mult_w_result_range320w(0) <= wire_man_product2_mult_result(5);
	wire_man_product2_mult_w_result_range323w(0) <= wire_man_product2_mult_result(6);
	wire_man_product2_mult_w_result_range326w(0) <= wire_man_product2_mult_result(7);
	wire_man_product2_mult_w_result_range329w(0) <= wire_man_product2_mult_result(8);
	wire_man_product2_mult_w_result_range332w(0) <= wire_man_product2_mult_result(9);
	man_product2_mult :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 24,
		LPM_WIDTHB => 24,
		LPM_WIDTHP => 48,
		LPM_WIDTHS => 1,
		lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES"
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_man_product2_mult_dataa,
		datab => wire_man_product2_mult_datab,
		result => wire_man_product2_mult_result
	  );

 END RTL; --fp_mult_altfp_mult_v9o
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fp_mult IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END fp_mult;


ARCHITECTURE RTL OF fp_mult IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT fp_mult_altfp_mult_v9o
	PORT (
			aclr	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	fp_mult_altfp_mult_v9o_component : fp_mult_altfp_mult_v9o
	PORT MAP (
		aclr => aclr,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: FPM_FORMAT STRING "Single"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "YES"
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: EXCEPTION_HANDLING STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_mult"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "5"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_mult.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
